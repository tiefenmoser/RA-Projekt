library ieee;
use ieee.std_logic_1164.all;


use work.Constant_Package.all;

entity alu is
    port(
        

    );
end alu;   


