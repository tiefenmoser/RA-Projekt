entity hello is
end entity hello;
architecture arc of hello is
begin
assert false report "Willkommen zu GdTI!" severity note;
end architecture arc;
