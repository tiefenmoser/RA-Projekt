library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constant_package.all;

entity sltu is
end sltu;



architecture behave of sltu is
    begin
end architecture;